desc_sv=AdFreeZone-loggning
