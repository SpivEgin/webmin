desc_sv=AdFreeZone-serverindex
